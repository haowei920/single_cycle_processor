import rv32i_types::*;
